`include "uvm_macros.svh"

package apbm_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  //`include "define.svh"
  `include "apbm_sequence_item.sv"
  `include "apbm_sequence.sv"
  `include "apbm_sequencer.sv"
  `include "apbm_driver.sv"
  `include "apbm_active_monitor.sv"
  `include "apbm_passive_monitor.sv"
  `include "apbm_active_agent.sv"
  `include "apbm_passive_agent.sv"
  `include "apbm_scoreboard.sv"
  //`include "apbm_subscriber.sv"
  `include "apbm_environment.sv"
  `include "apbm_test.sv"
endpackage
